module commit(
    );
